-- testRam_GN.vhd

-- Generated using ACDS version 16.0 222

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity testRam_GN is
	port (
		Avalon_ST_Source_ready         : in  std_logic                     := '0';             --         Avalon_ST_Source_ready.wire
		Clock                          : in  std_logic                     := '0';             --                          Clock.clk
		aclr                           : in  std_logic                     := '0';             --                               .reset_n
		Input                          : in  std_logic_vector(17 downto 0) := (others => '0'); --                          Input.wire
		Avalon_ST_Sink_endofpacket     : in  std_logic                     := '0';             --     Avalon_ST_Sink_endofpacket.wire
		Avalon_ST_Source_endofpacket   : out std_logic;                                        --   Avalon_ST_Source_endofpacket.wire
		Avalon_ST_Sink_ready           : out std_logic;                                        --           Avalon_ST_Sink_ready.wire
		Avalon_ST_Source_valid         : out std_logic;                                        --         Avalon_ST_Source_valid.wire
		Avalon_ST_Sink_data            : in  std_logic_vector(23 downto 0) := (others => '0'); --            Avalon_ST_Sink_data.wire
		Avalon_ST_Source_data          : out std_logic_vector(23 downto 0);                    --          Avalon_ST_Source_data.wire
		Avalon_ST_Sink_startofpacket   : in  std_logic                     := '0';             --   Avalon_ST_Sink_startofpacket.wire
		Avalon_ST_Sink_valid           : in  std_logic                     := '0';             --           Avalon_ST_Sink_valid.wire
		Avalon_ST_Source_startofpacket : out std_logic                                         -- Avalon_ST_Source_startofpacket.wire
	);
end entity testRam_GN;

architecture rtl of testRam_GN is
	component alt_dspbuilder_clock_GNF343OQUJ is
		port (
			aclr      : in  std_logic := 'X'; -- reset
			aclr_n    : in  std_logic := 'X'; -- reset_n
			aclr_out  : out std_logic;        -- reset
			clock     : in  std_logic := 'X'; -- clk
			clock_out : out std_logic         -- clk
		);
	end component alt_dspbuilder_clock_GNF343OQUJ;

	component alt_dspbuilder_port_GN37ALZBS4 is
		port (
			input  : in  std_logic := 'X'; -- wire
			output : out std_logic         -- wire
		);
	end component alt_dspbuilder_port_GN37ALZBS4;

	component alt_dspbuilder_port_GNOC3SGKQJ is
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(23 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNOC3SGKQJ;

	component alt_dspbuilder_port_GN2CABCRLL is
		port (
			input  : in  std_logic_vector(17 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(17 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GN2CABCRLL;

	component testRam_GN_testRam_ram is
		port (
			valid_in  : in  std_logic                     := 'X';             -- wire
			valid_out : out std_logic;                                        -- wire
			sof_in    : in  std_logic                     := 'X';             -- wire
			eof_in    : in  std_logic                     := 'X';             -- wire
			eof_out   : out std_logic_vector(0 downto 0);                     -- wire
			sof_out   : out std_logic_vector(0 downto 0);                     -- wire
			Clock     : in  std_logic                     := 'X';             -- clk
			aclr      : in  std_logic                     := 'X';             -- reset
			pixel_in  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			control   : in  std_logic_vector(17 downto 0) := (others => 'X'); -- wire
			pixel_out : out std_logic_vector(23 downto 0)                     -- wire
		);
	end component testRam_GN_testRam_ram;

	component alt_dspbuilder_cast_GNSB3OXIQS is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(0 downto 0) := (others => 'X'); -- wire
			output : out std_logic                                        -- wire
		);
	end component alt_dspbuilder_cast_GNSB3OXIQS;

	signal avalon_st_source_ready_0_output_wire       : std_logic;                     -- Avalon_ST_Source_ready_0:output -> Avalon_ST_Sink_ready_0:input
	signal avalon_st_sink_data_0_output_wire          : std_logic_vector(23 downto 0); -- Avalon_ST_Sink_data_0:output -> testRam_ram_0:pixel_in
	signal avalon_st_sink_valid_0_output_wire         : std_logic;                     -- Avalon_ST_Sink_valid_0:output -> testRam_ram_0:valid_in
	signal avalon_st_sink_startofpacket_0_output_wire : std_logic;                     -- Avalon_ST_Sink_startofpacket_0:output -> testRam_ram_0:sof_in
	signal avalon_st_sink_endofpacket_0_output_wire   : std_logic;                     -- Avalon_ST_Sink_endofpacket_0:output -> testRam_ram_0:eof_in
	signal input_0_output_wire                        : std_logic_vector(17 downto 0); -- Input_0:output -> testRam_ram_0:control
	signal testram_ram_0_pixel_out_wire               : std_logic_vector(23 downto 0); -- testRam_ram_0:pixel_out -> Avalon_ST_Source_data_0:input
	signal testram_ram_0_valid_out_wire               : std_logic;                     -- testRam_ram_0:valid_out -> Avalon_ST_Source_valid_0:input
	signal testram_ram_0_sof_out_wire                 : std_logic_vector(0 downto 0);  -- testRam_ram_0:sof_out -> cast5:input
	signal cast5_output_wire                          : std_logic;                     -- cast5:output -> Avalon_ST_Source_startofpacket_0:input
	signal testram_ram_0_eof_out_wire                 : std_logic_vector(0 downto 0);  -- testRam_ram_0:eof_out -> cast6:input
	signal cast6_output_wire                          : std_logic;                     -- cast6:output -> Avalon_ST_Source_endofpacket_0:input
	signal clock_0_clock_output_clk                   : std_logic;                     -- Clock_0:clock_out -> testRam_ram_0:Clock
	signal clock_0_clock_output_reset                 : std_logic;                     -- Clock_0:aclr_out -> testRam_ram_0:aclr

begin

	clock_0 : component alt_dspbuilder_clock_GNF343OQUJ
		port map (
			clock_out => clock_0_clock_output_clk,   -- clock_output.clk
			aclr_out  => clock_0_clock_output_reset, --             .reset
			clock     => Clock,                      --        clock.clk
			aclr_n    => aclr                        --             .reset_n
		);

	avalon_st_sink_valid_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => Avalon_ST_Sink_valid,               --  input.wire
			output => avalon_st_sink_valid_0_output_wire  -- output.wire
		);

	avalon_st_source_data_0 : component alt_dspbuilder_port_GNOC3SGKQJ
		port map (
			input  => testram_ram_0_pixel_out_wire, --  input.wire
			output => Avalon_ST_Source_data         -- output.wire
		);

	avalon_st_sink_endofpacket_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => Avalon_ST_Sink_endofpacket,               --  input.wire
			output => avalon_st_sink_endofpacket_0_output_wire  -- output.wire
		);

	avalon_st_source_ready_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => Avalon_ST_Source_ready,               --  input.wire
			output => avalon_st_source_ready_0_output_wire  -- output.wire
		);

	input_0 : component alt_dspbuilder_port_GN2CABCRLL
		port map (
			input  => Input,               --  input.wire
			output => input_0_output_wire  -- output.wire
		);

	testram_ram_0 : component testRam_GN_testRam_ram
		port map (
			valid_in  => avalon_st_sink_valid_0_output_wire,         --  valid_in.wire
			valid_out => testram_ram_0_valid_out_wire,               -- valid_out.wire
			sof_in    => avalon_st_sink_startofpacket_0_output_wire, --    sof_in.wire
			eof_in    => avalon_st_sink_endofpacket_0_output_wire,   --    eof_in.wire
			eof_out   => testram_ram_0_eof_out_wire,                 --   eof_out.wire
			sof_out   => testram_ram_0_sof_out_wire,                 --   sof_out.wire
			Clock     => clock_0_clock_output_clk,                   --     Clock.clk
			aclr      => clock_0_clock_output_reset,                 --          .reset
			pixel_in  => avalon_st_sink_data_0_output_wire,          --  pixel_in.wire
			control   => input_0_output_wire,                        --   control.wire
			pixel_out => testram_ram_0_pixel_out_wire                -- pixel_out.wire
		);

	avalon_st_source_endofpacket_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => cast6_output_wire,            --  input.wire
			output => Avalon_ST_Source_endofpacket  -- output.wire
		);

	avalon_st_sink_startofpacket_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => Avalon_ST_Sink_startofpacket,               --  input.wire
			output => avalon_st_sink_startofpacket_0_output_wire  -- output.wire
		);

	avalon_st_source_valid_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => testram_ram_0_valid_out_wire, --  input.wire
			output => Avalon_ST_Source_valid        -- output.wire
		);

	avalon_st_sink_data_0 : component alt_dspbuilder_port_GNOC3SGKQJ
		port map (
			input  => Avalon_ST_Sink_data,               --  input.wire
			output => avalon_st_sink_data_0_output_wire  -- output.wire
		);

	avalon_st_sink_ready_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => avalon_st_source_ready_0_output_wire, --  input.wire
			output => Avalon_ST_Sink_ready                  -- output.wire
		);

	avalon_st_source_startofpacket_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => cast5_output_wire,              --  input.wire
			output => Avalon_ST_Source_startofpacket  -- output.wire
		);

	cast5 : component alt_dspbuilder_cast_GNSB3OXIQS
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => testram_ram_0_sof_out_wire, --  input.wire
			output => cast5_output_wire           -- output.wire
		);

	cast6 : component alt_dspbuilder_cast_GNSB3OXIQS
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => testram_ram_0_eof_out_wire, --  input.wire
			output => cast6_output_wire           -- output.wire
		);

end architecture rtl; -- of testRam_GN
