-- testRam_GN_testRam_ram.vhd

-- Generated using ACDS version 16.0 222

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity testRam_GN_testRam_ram is
	port (
		valid_in  : in  std_logic                     := '0';             --  valid_in.wire
		valid_out : out std_logic;                                        -- valid_out.wire
		sof_in    : in  std_logic                     := '0';             --    sof_in.wire
		eof_in    : in  std_logic                     := '0';             --    eof_in.wire
		eof_out   : out std_logic_vector(0 downto 0);                     --   eof_out.wire
		sof_out   : out std_logic_vector(0 downto 0);                     --   sof_out.wire
		Clock     : in  std_logic                     := '0';             --     Clock.clk
		aclr      : in  std_logic                     := '0';             --          .reset
		pixel_in  : in  std_logic_vector(23 downto 0) := (others => '0'); --  pixel_in.wire
		control   : in  std_logic_vector(17 downto 0) := (others => '0'); --   control.wire
		pixel_out : out std_logic_vector(23 downto 0)                     -- pixel_out.wire
	);
end entity testRam_GN_testRam_ram;

architecture rtl of testRam_GN_testRam_ram is
	component alt_dspbuilder_clock_GNQFU4PUDH is
		port (
			aclr      : in  std_logic := 'X'; -- reset
			aclr_n    : in  std_logic := 'X'; -- reset_n
			aclr_out  : out std_logic;        -- reset
			clock     : in  std_logic := 'X'; -- clk
			clock_out : out std_logic         -- clk
		);
	end component alt_dspbuilder_clock_GNQFU4PUDH;

	component alt_dspbuilder_port_GN37ALZBS4 is
		port (
			input  : in  std_logic := 'X'; -- wire
			output : out std_logic         -- wire
		);
	end component alt_dspbuilder_port_GN37ALZBS4;

	component alt_dspbuilder_port_GNXAOKDYKC is
		port (
			input  : in  std_logic_vector(0 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(0 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNXAOKDYKC;

	component alt_dspbuilder_multiplexer_GNAIWAHV3K is
		generic (
			number_inputs          : natural  := 4;
			pipeline               : natural  := 0;
			width                  : positive := 8;
			HDLTYPE                : string   := "STD_LOGIC_VECTOR";
			use_one_hot_select_bus : natural  := 0
		);
		port (
			clock     : in  std_logic                    := 'X';             -- clk
			aclr      : in  std_logic                    := 'X';             -- reset
			sel       : in  std_logic_vector(0 downto 0) := (others => 'X'); -- wire
			result    : out std_logic_vector(0 downto 0);                    -- wire
			ena       : in  std_logic                    := 'X';             -- wire
			user_aclr : in  std_logic                    := 'X';             -- wire
			in0       : in  std_logic_vector(0 downto 0) := (others => 'X'); -- wire
			in1       : in  std_logic_vector(0 downto 0) := (others => 'X')  -- wire
		);
	end component alt_dspbuilder_multiplexer_GNAIWAHV3K;

	component alt_dspbuilder_gnd_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_gnd_GN;

	component alt_dspbuilder_vcc_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_vcc_GN;

	component alt_dspbuilder_port_GNOC3SGKQJ is
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(23 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNOC3SGKQJ;

	component alt_dspbuilder_multiplexer_GNCALBUTDR is
		generic (
			number_inputs          : natural  := 4;
			pipeline               : natural  := 0;
			width                  : positive := 8;
			HDLTYPE                : string   := "STD_LOGIC_VECTOR";
			use_one_hot_select_bus : natural  := 0
		);
		port (
			clock     : in  std_logic                     := 'X';             -- clk
			aclr      : in  std_logic                     := 'X';             -- reset
			sel       : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- wire
			result    : out std_logic_vector(23 downto 0);                    -- wire
			ena       : in  std_logic                     := 'X';             -- wire
			user_aclr : in  std_logic                     := 'X';             -- wire
			in0       : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			in1       : in  std_logic_vector(23 downto 0) := (others => 'X')  -- wire
		);
	end component alt_dspbuilder_multiplexer_GNCALBUTDR;

	component alt_dspbuilder_delay_GNLRSWL7NV is
		generic (
			ClockPhase : string   := "1";
			BitPattern : string   := "00000001";
			width      : positive := 8;
			use_init   : natural  := 0;
			delay      : positive := 1
		);
		port (
			aclr   : in  std_logic                          := 'X';             -- clk
			clock  : in  std_logic                          := 'X';             -- clk
			ena    : in  std_logic                          := 'X';             -- wire
			input  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(width-1 downto 0);                    -- wire
			sclr   : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_delay_GNLRSWL7NV;

	component testRam_GN_testRam_ram_counter1 is
		port (
			Clock    : in  std_logic                     := 'X'; -- clk
			aclr     : in  std_logic                     := 'X'; -- reset
			valid_in : in  std_logic                     := 'X'; -- wire
			eof_in   : in  std_logic                     := 'X'; -- wire
			col_out  : out std_logic_vector(13 downto 0)         -- wire
		);
	end component testRam_GN_testRam_ram_counter1;

	component alt_dspbuilder_cast_GNA7YF6ZOH is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(17 downto 0) := (others => 'X'); -- wire
			output : out std_logic                                         -- wire
		);
	end component alt_dspbuilder_cast_GNA7YF6ZOH;

	component alt_dspbuilder_dualram_GNPI5EKKTA is
		generic (
			ClockPhase       : string   := "1";
			numwords         : positive := 3;
			register_outputs : natural  := 1;
			data_width       : positive := 8;
			supportROM       : natural  := 1;
			ram_block_type   : string   := "AUTO";
			use_ena          : natural  := 0;
			XFILE            : string   := "input.hex";
			initialization   : string   := "Blank";
			dont_care        : natural  := 0;
			family           : string   := "STRATIXV"
		);
		port (
			clock   : in  std_logic                     := 'X';             -- clk
			aclr    : in  std_logic                     := 'X';             -- reset
			data    : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			rd_addr : in  std_logic_vector(13 downto 0) := (others => 'X'); -- wire
			wr_addr : in  std_logic_vector(13 downto 0) := (others => 'X'); -- wire
			wren    : in  std_logic                     := 'X';             -- wire
			ena     : in  std_logic                     := 'X';             -- wire
			q       : out std_logic_vector(23 downto 0)                     -- wire
		);
	end component alt_dspbuilder_dualram_GNPI5EKKTA;

	component alt_dspbuilder_logical_bus_op_GNOC3X2UWP is
		generic (
			logical_op       : string   := "AltAND";
			lpm_width        : positive := 8;
			shift_amount     : natural  := 3;
			mask_value       : string   := "10101010";
			signextendrshift : natural  := 1
		);
		port (
			dataa  : in  std_logic_vector(lpm_width-1 downto 0) := (others => 'X'); -- wire
			result : out std_logic_vector(lpm_width-1 downto 0)                     -- wire
		);
	end component alt_dspbuilder_logical_bus_op_GNOC3X2UWP;

	component alt_dspbuilder_delay_GNQBXYU75H is
		generic (
			ClockPhase : string   := "1";
			BitPattern : string   := "00000001";
			width      : positive := 8;
			use_init   : natural  := 0;
			delay      : positive := 1
		);
		port (
			aclr   : in  std_logic                          := 'X';             -- clk
			clock  : in  std_logic                          := 'X';             -- clk
			ena    : in  std_logic                          := 'X';             -- wire
			input  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(width-1 downto 0);                    -- wire
			sclr   : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_delay_GNQBXYU75H;

	component alt_dspbuilder_port_GN2CABCRLL is
		port (
			input  : in  std_logic_vector(17 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(17 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GN2CABCRLL;

	component testRam_GN_testRam_ram_counter is
		port (
			valid_in : in  std_logic                     := 'X'; -- wire
			eof_in   : in  std_logic                     := 'X'; -- wire
			col_out  : out std_logic_vector(13 downto 0);        -- wire
			Clock    : in  std_logic                     := 'X'; -- clk
			aclr     : in  std_logic                     := 'X'  -- reset
		);
	end component testRam_GN_testRam_ram_counter;

	component alt_dspbuilder_dualram_GNYFEXMTMW is
		generic (
			ClockPhase       : string   := "1";
			numwords         : positive := 3;
			register_outputs : natural  := 1;
			data_width       : positive := 8;
			supportROM       : natural  := 1;
			ram_block_type   : string   := "AUTO";
			use_ena          : natural  := 0;
			XFILE            : string   := "input.hex";
			initialization   : string   := "Blank";
			dont_care        : natural  := 0;
			family           : string   := "STRATIXV"
		);
		port (
			clock   : in  std_logic                     := 'X';             -- clk
			aclr    : in  std_logic                     := 'X';             -- reset
			data    : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			rd_addr : in  std_logic_vector(13 downto 0) := (others => 'X'); -- wire
			wr_addr : in  std_logic_vector(13 downto 0) := (others => 'X'); -- wire
			wren    : in  std_logic                     := 'X';             -- wire
			ena     : in  std_logic                     := 'X';             -- wire
			q       : out std_logic_vector(23 downto 0)                     -- wire
		);
	end component alt_dspbuilder_dualram_GNYFEXMTMW;

	component alt_dspbuilder_delay_GNGQ56ZS4N is
		generic (
			ClockPhase : string   := "1";
			BitPattern : string   := "00000001";
			width      : positive := 8;
			use_init   : natural  := 0;
			delay      : positive := 1
		);
		port (
			aclr   : in  std_logic                          := 'X';             -- clk
			clock  : in  std_logic                          := 'X';             -- clk
			ena    : in  std_logic                          := 'X';             -- wire
			input  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(width-1 downto 0);                    -- wire
			sclr   : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_delay_GNGQ56ZS4N;

	component alt_dspbuilder_cast_GN46N4UJ5S is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic                    := 'X'; -- wire
			output : out std_logic_vector(0 downto 0)         -- wire
		);
	end component alt_dspbuilder_cast_GN46N4UJ5S;

	signal multiplexeruser_aclrgnd_output_wire  : std_logic;                     -- Multiplexeruser_aclrGND:output -> Multiplexer:user_aclr
	signal multiplexerenavcc_output_wire        : std_logic;                     -- MultiplexerenaVCC:output -> Multiplexer:ena
	signal multiplexer1user_aclrgnd_output_wire : std_logic;                     -- Multiplexer1user_aclrGND:output -> Multiplexer1:user_aclr
	signal multiplexer1enavcc_output_wire       : std_logic;                     -- Multiplexer1enaVCC:output -> Multiplexer1:ena
	signal multiplexer2user_aclrgnd_output_wire : std_logic;                     -- Multiplexer2user_aclrGND:output -> Multiplexer2:user_aclr
	signal multiplexer2enavcc_output_wire       : std_logic;                     -- Multiplexer2enaVCC:output -> Multiplexer2:ena
	signal delaysclrgnd_output_wire             : std_logic;                     -- DelaysclrGND:output -> Delay:sclr
	signal dual_port_ram1enavcc_output_wire     : std_logic;                     -- Dual_Port_RAM1enaVCC:output -> Dual_Port_RAM1:ena
	signal delay2sclrgnd_output_wire            : std_logic;                     -- Delay2sclrGND:output -> Delay2:sclr
	signal delay1sclrgnd_output_wire            : std_logic;                     -- Delay1sclrGND:output -> Delay1:sclr
	signal dual_port_ramenavcc_output_wire      : std_logic;                     -- Dual_Port_RAMenaVCC:output -> Dual_Port_RAM:ena
	signal delay5sclrgnd_output_wire            : std_logic;                     -- Delay5sclrGND:output -> Delay5:sclr
	signal delay4sclrgnd_output_wire            : std_logic;                     -- Delay4sclrGND:output -> Delay4:sclr
	signal delay3sclrgnd_output_wire            : std_logic;                     -- Delay3sclrGND:output -> Delay3:sclr
	signal delay1_output_wire                   : std_logic_vector(0 downto 0);  -- Delay1:output -> [Delay3:input, Multiplexer:in0]
	signal delay4_output_wire                   : std_logic_vector(0 downto 0);  -- Delay4:output -> [Delay5:input, Multiplexer1:in0]
	signal delay_output_wire                    : std_logic_vector(13 downto 0); -- Delay:output -> Dual_Port_RAM:wr_addr
	signal delay2_output_wire                   : std_logic_vector(13 downto 0); -- Delay2:output -> Dual_Port_RAM1:wr_addr
	signal testram_ram_counter_0_col_out_wire   : std_logic_vector(13 downto 0); -- testRam_ram_counter_0:col_out -> [Dual_Port_RAM1:rd_addr, Dual_Port_RAM:rd_addr]
	signal pixel_in_0_output_wire               : std_logic_vector(23 downto 0); -- pixel_in_0:output -> [Dual_Port_RAM1:data, Dual_Port_RAM:data]
	signal valid_in_0_output_wire               : std_logic;                     -- valid_in_0:output -> [Delay1:ena, Delay2:ena, Delay3:ena, Delay4:ena, Delay5:ena, Delay:ena, Dual_Port_RAM1:wren, Dual_Port_RAM:wren, testRam_ram_counter1_0:valid_in, testRam_ram_counter_0:valid_in, valid_out_0:input]
	signal control_0_output_wire                : std_logic_vector(17 downto 0); -- control_0:output -> [AltBus1:input, AltBus:input, Logical_Bus_Operator:dataa]
	signal testram_ram_counter1_0_col_out_wire  : std_logic_vector(13 downto 0); -- testRam_ram_counter1_0:col_out -> [Delay2:input, Delay:input]
	signal logical_bus_operator_result_wire     : std_logic_vector(17 downto 0); -- Logical_Bus_Operator:result -> AltBus2:input
	signal delay3_output_wire                   : std_logic_vector(0 downto 0);  -- Delay3:output -> Multiplexer:in1
	signal delay5_output_wire                   : std_logic_vector(0 downto 0);  -- Delay5:output -> Multiplexer1:in1
	signal dual_port_ram1_q_wire                : std_logic_vector(23 downto 0); -- Dual_Port_RAM1:q -> Multiplexer2:in0
	signal dual_port_ram_q_wire                 : std_logic_vector(23 downto 0); -- Dual_Port_RAM:q -> Multiplexer2:in1
	signal eof_in_0_output_wire                 : std_logic;                     -- eof_in_0:output -> [cast1:input, testRam_ram_counter1_0:eof_in, testRam_ram_counter_0:eof_in]
	signal multiplexer2_result_wire             : std_logic_vector(23 downto 0); -- Multiplexer2:result -> pixel_out_0:input
	signal multiplexer1_result_wire             : std_logic_vector(0 downto 0);  -- Multiplexer1:result -> sof_out_0:input
	signal multiplexer_result_wire              : std_logic_vector(0 downto 0);  -- Multiplexer:result -> eof_out_0:input
	signal sof_in_0_output_wire                 : std_logic;                     -- sof_in_0:output -> cast0:input
	signal cast0_output_wire                    : std_logic_vector(0 downto 0);  -- cast0:output -> Delay4:input
	signal cast1_output_wire                    : std_logic_vector(0 downto 0);  -- cast1:output -> Delay1:input
	signal altbus_output_wire                   : std_logic;                     -- AltBus:output -> cast2:input
	signal cast2_output_wire                    : std_logic_vector(0 downto 0);  -- cast2:output -> Multiplexer:sel
	signal altbus1_output_wire                  : std_logic;                     -- AltBus1:output -> cast3:input
	signal cast3_output_wire                    : std_logic_vector(0 downto 0);  -- cast3:output -> Multiplexer1:sel
	signal altbus2_output_wire                  : std_logic;                     -- AltBus2:output -> cast4:input
	signal cast4_output_wire                    : std_logic_vector(0 downto 0);  -- cast4:output -> Multiplexer2:sel
	signal clock_0_clock_output_clk             : std_logic;                     -- Clock_0:clock_out -> [Delay1:clock, Delay2:clock, Delay3:clock, Delay4:clock, Delay5:clock, Delay:clock, Dual_Port_RAM1:clock, Dual_Port_RAM:clock, Multiplexer1:clock, Multiplexer2:clock, Multiplexer:clock, testRam_ram_counter1_0:Clock, testRam_ram_counter_0:Clock]
	signal clock_0_clock_output_reset           : std_logic;                     -- Clock_0:aclr_out -> [Delay1:aclr, Delay2:aclr, Delay3:aclr, Delay4:aclr, Delay5:aclr, Delay:aclr, Dual_Port_RAM1:aclr, Dual_Port_RAM:aclr, Multiplexer1:aclr, Multiplexer2:aclr, Multiplexer:aclr, testRam_ram_counter1_0:aclr, testRam_ram_counter_0:aclr]

begin

	clock_0 : component alt_dspbuilder_clock_GNQFU4PUDH
		port map (
			clock_out => clock_0_clock_output_clk,   -- clock_output.clk
			aclr_out  => clock_0_clock_output_reset, --             .reset
			clock     => Clock,                      --        clock.clk
			aclr      => aclr                        --             .reset
		);

	valid_in_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => valid_in,               --  input.wire
			output => valid_in_0_output_wire  -- output.wire
		);

	eof_out_0 : component alt_dspbuilder_port_GNXAOKDYKC
		port map (
			input  => multiplexer_result_wire, --  input.wire
			output => eof_out                  -- output.wire
		);

	multiplexer : component alt_dspbuilder_multiplexer_GNAIWAHV3K
		generic map (
			number_inputs          => 2,
			pipeline               => 0,
			width                  => 1,
			HDLTYPE                => "STD_LOGIC_VECTOR",
			use_one_hot_select_bus => 0
		)
		port map (
			clock     => clock_0_clock_output_clk,            -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,          --           .reset
			sel       => cast2_output_wire,                   --        sel.wire
			result    => multiplexer_result_wire,             --     result.wire
			ena       => multiplexerenavcc_output_wire,       --        ena.wire
			user_aclr => multiplexeruser_aclrgnd_output_wire, --  user_aclr.wire
			in0       => delay1_output_wire,                  --        in0.wire
			in1       => delay3_output_wire                   --        in1.wire
		);

	multiplexeruser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplexeruser_aclrgnd_output_wire  -- output.wire
		);

	multiplexerenavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplexerenavcc_output_wire  -- output.wire
		);

	multiplexer1 : component alt_dspbuilder_multiplexer_GNAIWAHV3K
		generic map (
			number_inputs          => 2,
			pipeline               => 0,
			width                  => 1,
			HDLTYPE                => "STD_LOGIC_VECTOR",
			use_one_hot_select_bus => 0
		)
		port map (
			clock     => clock_0_clock_output_clk,             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,           --           .reset
			sel       => cast3_output_wire,                    --        sel.wire
			result    => multiplexer1_result_wire,             --     result.wire
			ena       => multiplexer1enavcc_output_wire,       --        ena.wire
			user_aclr => multiplexer1user_aclrgnd_output_wire, --  user_aclr.wire
			in0       => delay4_output_wire,                   --        in0.wire
			in1       => delay5_output_wire                    --        in1.wire
		);

	multiplexer1user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplexer1user_aclrgnd_output_wire  -- output.wire
		);

	multiplexer1enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplexer1enavcc_output_wire  -- output.wire
		);

	pixel_in_0 : component alt_dspbuilder_port_GNOC3SGKQJ
		port map (
			input  => pixel_in,               --  input.wire
			output => pixel_in_0_output_wire  -- output.wire
		);

	multiplexer2 : component alt_dspbuilder_multiplexer_GNCALBUTDR
		generic map (
			number_inputs          => 2,
			pipeline               => 0,
			width                  => 24,
			HDLTYPE                => "STD_LOGIC_VECTOR",
			use_one_hot_select_bus => 0
		)
		port map (
			clock     => clock_0_clock_output_clk,             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,           --           .reset
			sel       => cast4_output_wire,                    --        sel.wire
			result    => multiplexer2_result_wire,             --     result.wire
			ena       => multiplexer2enavcc_output_wire,       --        ena.wire
			user_aclr => multiplexer2user_aclrgnd_output_wire, --  user_aclr.wire
			in0       => dual_port_ram1_q_wire,                --        in0.wire
			in1       => dual_port_ram_q_wire                  --        in1.wire
		);

	multiplexer2user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplexer2user_aclrgnd_output_wire  -- output.wire
		);

	multiplexer2enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplexer2enavcc_output_wire  -- output.wire
		);

	delay : component alt_dspbuilder_delay_GNLRSWL7NV
		generic map (
			ClockPhase => "1",
			BitPattern => "00000000000001",
			width      => 14,
			use_init   => 0,
			delay      => 2
		)
		port map (
			input  => testram_ram_counter1_0_col_out_wire, --      input.wire
			clock  => clock_0_clock_output_clk,            -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,          --           .reset
			output => delay_output_wire,                   --     output.wire
			sclr   => delaysclrgnd_output_wire,            --       sclr.wire
			ena    => valid_in_0_output_wire               --        ena.wire
		);

	delaysclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delaysclrgnd_output_wire  -- output.wire
		);

	valid_out_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => valid_in_0_output_wire, --  input.wire
			output => valid_out               -- output.wire
		);

	testram_ram_counter1_0 : component testRam_GN_testRam_ram_counter1
		port map (
			Clock    => clock_0_clock_output_clk,            --    Clock.clk
			aclr     => clock_0_clock_output_reset,          --         .reset
			valid_in => valid_in_0_output_wire,              -- valid_in.wire
			eof_in   => eof_in_0_output_wire,                --   eof_in.wire
			col_out  => testram_ram_counter1_0_col_out_wire  --  col_out.wire
		);

	altbus1 : component alt_dspbuilder_cast_GNA7YF6ZOH
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => control_0_output_wire, --  input.wire
			output => altbus1_output_wire    -- output.wire
		);

	dual_port_ram1 : component alt_dspbuilder_dualram_GNPI5EKKTA
		generic map (
			ClockPhase       => "1",
			numwords         => 10000,
			register_outputs => 1,
			data_width       => 24,
			supportROM       => 1,
			ram_block_type   => "M10K",
			use_ena          => 0,
			XFILE            => "input.hex",
			initialization   => "Blank",
			dont_care        => 1,
			family           => "Cyclone IV GX"
		)
		port map (
			clock   => clock_0_clock_output_clk,           -- clock_aclr.clk
			aclr    => clock_0_clock_output_reset,         --           .reset
			data    => pixel_in_0_output_wire,             --       data.wire
			rd_addr => testram_ram_counter_0_col_out_wire, --    rd_addr.wire
			wr_addr => delay2_output_wire,                 --    wr_addr.wire
			wren    => valid_in_0_output_wire,             --       wren.wire
			ena     => dual_port_ram1enavcc_output_wire,   --        ena.wire
			q       => dual_port_ram1_q_wire               --          q.wire
		);

	dual_port_ram1enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => dual_port_ram1enavcc_output_wire  -- output.wire
		);

	altbus2 : component alt_dspbuilder_cast_GNA7YF6ZOH
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => logical_bus_operator_result_wire, --  input.wire
			output => altbus2_output_wire               -- output.wire
		);

	logical_bus_operator : component alt_dspbuilder_logical_bus_op_GNOC3X2UWP
		generic map (
			logical_op       => "AltShiftRight",
			lpm_width        => 18,
			shift_amount     => 1,
			mask_value       => "111111111111111011",
			signextendrshift => 0
		)
		port map (
			dataa  => control_0_output_wire,            --  dataa.wire
			result => logical_bus_operator_result_wire  -- result.wire
		);

	delay2 : component alt_dspbuilder_delay_GNLRSWL7NV
		generic map (
			ClockPhase => "1",
			BitPattern => "00000000000001",
			width      => 14,
			use_init   => 0,
			delay      => 2
		)
		port map (
			input  => testram_ram_counter1_0_col_out_wire, --      input.wire
			clock  => clock_0_clock_output_clk,            -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,          --           .reset
			output => delay2_output_wire,                  --     output.wire
			sclr   => delay2sclrgnd_output_wire,           --       sclr.wire
			ena    => valid_in_0_output_wire               --        ena.wire
		);

	delay2sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay2sclrgnd_output_wire  -- output.wire
		);

	altbus : component alt_dspbuilder_cast_GNA7YF6ZOH
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => control_0_output_wire, --  input.wire
			output => altbus_output_wire     -- output.wire
		);

	delay1 : component alt_dspbuilder_delay_GNQBXYU75H
		generic map (
			ClockPhase => "1",
			BitPattern => "1",
			width      => 1,
			use_init   => 0,
			delay      => 4
		)
		port map (
			input  => cast1_output_wire,          --      input.wire
			clock  => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset, --           .reset
			output => delay1_output_wire,         --     output.wire
			sclr   => delay1sclrgnd_output_wire,  --       sclr.wire
			ena    => valid_in_0_output_wire      --        ena.wire
		);

	delay1sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay1sclrgnd_output_wire  -- output.wire
		);

	control_0 : component alt_dspbuilder_port_GN2CABCRLL
		port map (
			input  => control,               --  input.wire
			output => control_0_output_wire  -- output.wire
		);

	eof_in_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => eof_in,               --  input.wire
			output => eof_in_0_output_wire  -- output.wire
		);

	testram_ram_counter_0 : component testRam_GN_testRam_ram_counter
		port map (
			valid_in => valid_in_0_output_wire,             -- valid_in.wire
			eof_in   => eof_in_0_output_wire,               --   eof_in.wire
			col_out  => testram_ram_counter_0_col_out_wire, --  col_out.wire
			Clock    => clock_0_clock_output_clk,           --    Clock.clk
			aclr     => clock_0_clock_output_reset          --         .reset
		);

	sof_in_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => sof_in,               --  input.wire
			output => sof_in_0_output_wire  -- output.wire
		);

	dual_port_ram : component alt_dspbuilder_dualram_GNYFEXMTMW
		generic map (
			ClockPhase       => "1",
			numwords         => 10000,
			register_outputs => 1,
			data_width       => 24,
			supportROM       => 1,
			ram_block_type   => "M10K",
			use_ena          => 0,
			XFILE            => "input.hex",
			initialization   => "Blank",
			dont_care        => 0,
			family           => "Cyclone IV GX"
		)
		port map (
			clock   => clock_0_clock_output_clk,           -- clock_aclr.clk
			aclr    => clock_0_clock_output_reset,         --           .reset
			data    => pixel_in_0_output_wire,             --       data.wire
			rd_addr => testram_ram_counter_0_col_out_wire, --    rd_addr.wire
			wr_addr => delay_output_wire,                  --    wr_addr.wire
			wren    => valid_in_0_output_wire,             --       wren.wire
			ena     => dual_port_ramenavcc_output_wire,    --        ena.wire
			q       => dual_port_ram_q_wire                --          q.wire
		);

	dual_port_ramenavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => dual_port_ramenavcc_output_wire  -- output.wire
		);

	delay5 : component alt_dspbuilder_delay_GNGQ56ZS4N
		generic map (
			ClockPhase => "1",
			BitPattern => "1",
			width      => 1,
			use_init   => 0,
			delay      => 1
		)
		port map (
			input  => delay4_output_wire,         --      input.wire
			clock  => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset, --           .reset
			output => delay5_output_wire,         --     output.wire
			sclr   => delay5sclrgnd_output_wire,  --       sclr.wire
			ena    => valid_in_0_output_wire      --        ena.wire
		);

	delay5sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay5sclrgnd_output_wire  -- output.wire
		);

	sof_out_0 : component alt_dspbuilder_port_GNXAOKDYKC
		port map (
			input  => multiplexer1_result_wire, --  input.wire
			output => sof_out                   -- output.wire
		);

	delay4 : component alt_dspbuilder_delay_GNQBXYU75H
		generic map (
			ClockPhase => "1",
			BitPattern => "1",
			width      => 1,
			use_init   => 0,
			delay      => 4
		)
		port map (
			input  => cast0_output_wire,          --      input.wire
			clock  => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset, --           .reset
			output => delay4_output_wire,         --     output.wire
			sclr   => delay4sclrgnd_output_wire,  --       sclr.wire
			ena    => valid_in_0_output_wire      --        ena.wire
		);

	delay4sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay4sclrgnd_output_wire  -- output.wire
		);

	pixel_out_0 : component alt_dspbuilder_port_GNOC3SGKQJ
		port map (
			input  => multiplexer2_result_wire, --  input.wire
			output => pixel_out                 -- output.wire
		);

	delay3 : component alt_dspbuilder_delay_GNGQ56ZS4N
		generic map (
			ClockPhase => "1",
			BitPattern => "1",
			width      => 1,
			use_init   => 0,
			delay      => 1
		)
		port map (
			input  => delay1_output_wire,         --      input.wire
			clock  => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset, --           .reset
			output => delay3_output_wire,         --     output.wire
			sclr   => delay3sclrgnd_output_wire,  --       sclr.wire
			ena    => valid_in_0_output_wire      --        ena.wire
		);

	delay3sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay3sclrgnd_output_wire  -- output.wire
		);

	cast0 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => sof_in_0_output_wire, --  input.wire
			output => cast0_output_wire     -- output.wire
		);

	cast1 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => eof_in_0_output_wire, --  input.wire
			output => cast1_output_wire     -- output.wire
		);

	cast2 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => altbus_output_wire, --  input.wire
			output => cast2_output_wire   -- output.wire
		);

	cast3 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => altbus1_output_wire, --  input.wire
			output => cast3_output_wire    -- output.wire
		);

	cast4 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => altbus2_output_wire, --  input.wire
			output => cast4_output_wire    -- output.wire
		);

end architecture rtl; -- of testRam_GN_testRam_ram
